`define N          8  
`define DATA_WIDTH 8
`define FIFO_DEPTH 8
parameter ADDR_WIDTH = $clog2(`FIFO_DEPTH);
                 
